module AND (y, a, b);

	input a, b;
	output y;

endmodule

module OR (y, a, b);

	input a, b;
	output y;

endmodule

module NOT (y, a);

	input a;
	output y;

endmodule

module DFF (CK, RS, D, Q);

	input CK, RS, D;
	output Q;

endmodule