module design1 (in1, in2, out1, out2);

	input in1, in2;
	output out1, out2;

	Test t1 (in1, in2, out1, out2);

endmodule