module top (a, c);

	input a, c;

endmodule
