module top (a, b, c, d);

	input a, b, c, d;
	
endmodule
	